$Generated from generate_tb.py
$
.include "/proj/cad/library/mosis/GF65_LPe/cmos10lpe_CDS_oa_dl064_11_20160415/models/YI-SM00030/Hspice/models/design.inc"

$.include dff.pex.sp $include your design
.option post runlvl=5

.param Tc=800p $CLK preiod 
.param Di=100p  $Input delay after rising edge of clock

$xi gnd! Q vdd! CLK R D design  $instantiate your design

vdd VDD! GND! 1.2v

vrst rst GND! PWL(0ps 0v 300ps 0v 350ps 1.2v 600ps 1.2v 650ps 0v) 
vclk clk GND! PULSE(0v 1.2v 0ps 50ps 50ps 'Tc/2-50ps' Tc)

$Expected Output:               D1:1011-D2:1011-   D3:-err-D4:0000-D5:0000-D6:0000-                    D7:1111-D8:-err-D9:0111-D10:1101
vin_ready in_ready GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' 0v 'Di+1*Tc' 0v 'Di+1*Tc+50ps' 0v 'Di+2*Tc' 0v 'Di+2*Tc+50ps' 1.2v 'Di+3*Tc' 1.2v 'Di+3*Tc+50ps' 0v 'Di+4*Tc' 0v 'Di+4*Tc+50ps' 0v 'Di+5*Tc' 0v 'Di+5*Tc+50ps' 0v 'Di+6*Tc' 0v 'Di+6*Tc+50ps' 0v 'Di+7*Tc' 0v 'Di+7*Tc+50ps' 0v 'Di+8*Tc' 0v 'Di+8*Tc+50ps' 0v 'Di+9*Tc' 0v 'Di+9*Tc+50ps' 0v 'Di+10*Tc' 0v 'Di+10*Tc+50ps' 1.2v 'Di+11*Tc' 1.2v 'Di+11*Tc+50ps' 0v 'Di+12*Tc' 0v 'Di+12*Tc+50ps' 0v 'Di+13*Tc' 0v 'Di+13*Tc+50ps' 0v 'Di+14*Tc' 0v 'Di+14*Tc+50ps' 0v 'Di+15*Tc' 0v 'Di+15*Tc+50ps' 0v 'Di+16*Tc' 0v 'Di+16*Tc+50ps' 0v 'Di+17*Tc' 0v 'Di+17*Tc+50ps' 0v 'Di+18*Tc' 0v 'Di+18*Tc+50ps' 0v 'Di+19*Tc' 0v 'Di+19*Tc+50ps' 0v 'Di+20*Tc' 0v 'Di+20*Tc+50ps' 0v 'Di+21*Tc' 0v 'Di+21*Tc+50ps' 1.2v 'Di+22*Tc' 1.2v 'Di+22*Tc+50ps' 0v 'Di+23*Tc' 0v 'Di+23*Tc+50ps' 0v 'Di+24*Tc' 0v 'Di+24*Tc+50ps' 0v 'Di+25*Tc' 0v 'Di+25*Tc+50ps' 0v 'Di+26*Tc' 0v 'Di+26*Tc+50ps' 0v 'Di+27*Tc' 0v 'Di+27*Tc+50ps' 0v 'Di+28*Tc' 0v 'Di+28*Tc+50ps' 0v 'Di+29*Tc' 0v 'Di+29*Tc+50ps' 1.2v 'Di+30*Tc' 1.2v 'Di+30*Tc+50ps' 0v 'Di+31*Tc' 0v 'Di+31*Tc+50ps' 0v 'Di+32*Tc' 0v 'Di+32*Tc+50ps' 0v 'Di+33*Tc' 0v 'Di+33*Tc+50ps' 0v 'Di+34*Tc' 0v 'Di+34*Tc+50ps' 0v 'Di+35*Tc' 0v 'Di+35*Tc+50ps' 0v 'Di+36*Tc' 0v 'Di+36*Tc+50ps' 0v 'Di+37*Tc' 0v 'Di+37*Tc+50ps' 1.2v 'Di+38*Tc' 1.2v 'Di+38*Tc+50ps' 0v 'Di+39*Tc' 0v 'Di+39*Tc+50ps' 0v 'Di+40*Tc' 0v 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' 0v 'Di+42*Tc' 0v 'Di+42*Tc+50ps' 0v 'Di+43*Tc' 0v 'Di+43*Tc+50ps' 0v 'Di+44*Tc' 0v 'Di+44*Tc+50ps' 0v 'Di+45*Tc' 0v 'Di+45*Tc+50ps' 1.2v 'Di+46*Tc' 1.2v 'Di+46*Tc+50ps' 0v 'Di+47*Tc' 0v 'Di+47*Tc+50ps' 0v 'Di+48*Tc' 0v 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' 0v 'Di+50*Tc' 0v 'Di+50*Tc+50ps' 0v 'Di+51*Tc' 0v 'Di+51*Tc+50ps' 0v 'Di+52*Tc' 0v 'Di+52*Tc+50ps' 0v 'Di+53*Tc' 0v 'Di+53*Tc+50ps' 0v 'Di+54*Tc' 0v 'Di+54*Tc+50ps' 0v 'Di+55*Tc' 0v 'Di+55*Tc+50ps' 0v 'Di+56*Tc' 0v 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' 0v 'Di+58*Tc' 0v 'Di+58*Tc+50ps' 0v 'Di+59*Tc' 0v 'Di+59*Tc+50ps' 0v 'Di+60*Tc' 0v 'Di+60*Tc+50ps' 0v 'Di+61*Tc' 0v 'Di+61*Tc+50ps' 0v 'Di+62*Tc' 0v 'Di+62*Tc+50ps' 0v 'Di+63*Tc' 0v 'Di+63*Tc+50ps' 0v 'Di+64*Tc' 0v 'Di+64*Tc+50ps' 0v 'Di+65*Tc' 0v 'Di+65*Tc+50ps' 0v 'Di+66*Tc' 0v 'Di+66*Tc+50ps' 0v 'Di+67*Tc' 0v 'Di+67*Tc+50ps' 0v 'Di+68*Tc' 0v 'Di+68*Tc+50ps' 0v 'Di+69*Tc' 0v 'Di+69*Tc+50ps' 0v 'Di+70*Tc' 0v 'Di+70*Tc+50ps' 0v 'Di+71*Tc' 0v 'Di+71*Tc+50ps' 0v 'Di+72*Tc' 0v 'Di+72*Tc+50ps' 0v 'Di+73*Tc' 0v 'Di+73*Tc+50ps' 1.2v 'Di+74*Tc' 1.2v 'Di+74*Tc+50ps' 0v 'Di+75*Tc' 0v 'Di+75*Tc+50ps' 0v 'Di+76*Tc' 0v 'Di+76*Tc+50ps' 0v 'Di+77*Tc' 0v 'Di+77*Tc+50ps' 0v 'Di+78*Tc' 0v 'Di+78*Tc+50ps' 0v 'Di+79*Tc' 0v 'Di+79*Tc+50ps' 0v 'Di+80*Tc' 0v 'Di+80*Tc+50ps' 0v 'Di+81*Tc' 0v 'Di+81*Tc+50ps' 1.2v 'Di+82*Tc' 1.2v 'Di+82*Tc+50ps' 0v 'Di+83*Tc' 0v 'Di+83*Tc+50ps' 0v 'Di+84*Tc' 0v 'Di+84*Tc+50ps' 0v 'Di+85*Tc' 0v 'Di+85*Tc+50ps' 0v 'Di+86*Tc' 0v 'Di+86*Tc+50ps' 0v 'Di+87*Tc' 0v 'Di+87*Tc+50ps' 0v 'Di+88*Tc' 0v 'Di+88*Tc+50ps' 0v 'Di+89*Tc' 0v 'Di+89*Tc+50ps' 1.2v 'Di+90*Tc' 1.2v 'Di+90*Tc+50ps' 0v 'Di+91*Tc' 0v 'Di+91*Tc+50ps' 0v 'Di+92*Tc' 0v 'Di+92*Tc+50ps' 0v 'Di+93*Tc' 0v 'Di+93*Tc+50ps' 0v 'Di+94*Tc' 0v 'Di+94*Tc+50ps' 0v 'Di+95*Tc' 0v 'Di+95*Tc+50ps' 0v 'Di+96*Tc' 0v 'Di+96*Tc+50ps' 0v 'Di+97*Tc' 0v 'Di+97*Tc+50ps' 1.2v 'Di+98*Tc' 1.2v 'Di+98*Tc+50ps' 0v 'Di+99*Tc' 0v 'Di+99*Tc+50ps' 0v 'Di+100*Tc' 0v 'Di+100*Tc+50ps' 0v 'Di+101*Tc' 0v 'Di+101*Tc+50ps' 0v 'Di+102*Tc' 0v 'Di+102*Tc+50ps' 0v 'Di+103*Tc' 0v 'Di+103*Tc+50ps' 0v 'Di+104*Tc' 0v 'Di+104*Tc+50ps' 0v 'Di+105*Tc' 0v 'Di+105*Tc+50ps' 0v 'Di+106*Tc' 0v 'Di+106*Tc+50ps' 0v 'Di+107*Tc' 0v 'Di+107*Tc+50ps' 0v 'Di+108*Tc' 0v 'Di+108*Tc+50ps' 0v 'Di+109*Tc' 0v 'Di+109*Tc+50ps' 0v 'Di+110*Tc' 0v)
vin in GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' 0v 'Di+1*Tc' 0v 'Di+1*Tc+50ps' 0v 'Di+2*Tc' 0v 'Di+2*Tc+50ps' 0v 'Di+3*Tc' 0v 'Di+3*Tc+50ps' 1.2v 'Di+4*Tc' 1.2v 'Di+4*Tc+50ps' 0v 'Di+5*Tc' 0v 'Di+5*Tc+50ps' 1.2v 'Di+6*Tc' 1.2v 'Di+6*Tc+50ps' 0v 'Di+7*Tc' 0v 'Di+7*Tc+50ps' 1.2v 'Di+8*Tc' 1.2v 'Di+8*Tc+50ps' 0v 'Di+9*Tc' 0v 'Di+9*Tc+50ps' 1.2v 'Di+10*Tc' 1.2v 'Di+10*Tc+50ps' 0v 'Di+11*Tc' 0v 'Di+11*Tc+50ps' 0v 'Di+12*Tc' 0v 'Di+12*Tc+50ps' 0v 'Di+13*Tc' 0v 'Di+13*Tc+50ps' 1.2v 'Di+14*Tc' 1.2v 'Di+14*Tc+50ps' 0v 'Di+15*Tc' 0v 'Di+15*Tc+50ps' 1.2v 'Di+16*Tc' 1.2v 'Di+16*Tc+50ps' 0v 'Di+17*Tc' 0v 'Di+17*Tc+50ps' 1.2v 'Di+18*Tc' 1.2v 'Di+18*Tc+50ps' 0v 'Di+19*Tc' 0v 'Di+19*Tc+50ps' 0v 'Di+20*Tc' 0v 'Di+20*Tc+50ps' 0v 'Di+21*Tc' 0v 'Di+21*Tc+50ps' 0v 'Di+22*Tc' 0v 'Di+22*Tc+50ps' 0v 'Di+23*Tc' 0v 'Di+23*Tc+50ps' 0v 'Di+24*Tc' 0v 'Di+24*Tc+50ps' 1.2v 'Di+25*Tc' 1.2v 'Di+25*Tc+50ps' 0v 'Di+26*Tc' 0v 'Di+26*Tc+50ps' 1.2v 'Di+27*Tc' 1.2v 'Di+27*Tc+50ps' 0v 'Di+28*Tc' 0v 'Di+28*Tc+50ps' 0v 'Di+29*Tc' 0v 'Di+29*Tc+50ps' 0v 'Di+30*Tc' 0v 'Di+30*Tc+50ps' 0v 'Di+31*Tc' 0v 'Di+31*Tc+50ps' 0v 'Di+32*Tc' 0v 'Di+32*Tc+50ps' 0v 'Di+33*Tc' 0v 'Di+33*Tc+50ps' 0v 'Di+34*Tc' 0v 'Di+34*Tc+50ps' 0v 'Di+35*Tc' 0v 'Di+35*Tc+50ps' 0v 'Di+36*Tc' 0v 'Di+36*Tc+50ps' 0v 'Di+37*Tc' 0v 'Di+37*Tc+50ps' 0v 'Di+38*Tc' 0v 'Di+38*Tc+50ps' 0v 'Di+39*Tc' 0v 'Di+39*Tc+50ps' 0v 'Di+40*Tc' 0v 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' 0v 'Di+42*Tc' 0v 'Di+42*Tc+50ps' 1.2v 'Di+43*Tc' 1.2v 'Di+43*Tc+50ps' 0v 'Di+44*Tc' 0v 'Di+44*Tc+50ps' 0v 'Di+45*Tc' 0v 'Di+45*Tc+50ps' 0v 'Di+46*Tc' 0v 'Di+46*Tc+50ps' 0v 'Di+47*Tc' 0v 'Di+47*Tc+50ps' 0v 'Di+48*Tc' 0v 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' 0v 'Di+50*Tc' 0v 'Di+50*Tc+50ps' 0v 'Di+51*Tc' 0v 'Di+51*Tc+50ps' 0v 'Di+52*Tc' 0v 'Di+52*Tc+50ps' 1.2v 'Di+53*Tc' 1.2v 'Di+53*Tc+50ps' 0v 'Di+54*Tc' 0v 'Di+54*Tc+50ps' 0v 'Di+55*Tc' 0v 'Di+55*Tc+50ps' 0v 'Di+56*Tc' 0v 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' 0v 'Di+58*Tc' 0v 'Di+58*Tc+50ps' 0v 'Di+59*Tc' 0v 'Di+59*Tc+50ps' 0v 'Di+60*Tc' 0v 'Di+60*Tc+50ps' 0v 'Di+61*Tc' 0v 'Di+61*Tc+50ps' 0v 'Di+62*Tc' 0v 'Di+62*Tc+50ps' 0v 'Di+63*Tc' 0v 'Di+63*Tc+50ps' 0v 'Di+64*Tc' 0v 'Di+64*Tc+50ps' 0v 'Di+65*Tc' 0v 'Di+65*Tc+50ps' 0v 'Di+66*Tc' 0v 'Di+66*Tc+50ps' 0v 'Di+67*Tc' 0v 'Di+67*Tc+50ps' 0v 'Di+68*Tc' 0v 'Di+68*Tc+50ps' 0v 'Di+69*Tc' 0v 'Di+69*Tc+50ps' 0v 'Di+70*Tc' 0v 'Di+70*Tc+50ps' 0v 'Di+71*Tc' 0v 'Di+71*Tc+50ps' 0v 'Di+72*Tc' 0v 'Di+72*Tc+50ps' 0v 'Di+73*Tc' 0v 'Di+73*Tc+50ps' 1.2v 'Di+74*Tc' 1.2v 'Di+74*Tc+50ps' 1.2v 'Di+75*Tc' 1.2v 'Di+75*Tc+50ps' 1.2v 'Di+76*Tc' 1.2v 'Di+76*Tc+50ps' 1.2v 'Di+77*Tc' 1.2v 'Di+77*Tc+50ps' 1.2v 'Di+78*Tc' 1.2v 'Di+78*Tc+50ps' 1.2v 'Di+79*Tc' 1.2v 'Di+79*Tc+50ps' 1.2v 'Di+80*Tc' 1.2v 'Di+80*Tc+50ps' 1.2v 'Di+81*Tc' 1.2v 'Di+81*Tc+50ps' 0v 'Di+82*Tc' 0v 'Di+82*Tc+50ps' 0v 'Di+83*Tc' 0v 'Di+83*Tc+50ps' 0v 'Di+84*Tc' 0v 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' 0v 'Di+86*Tc' 0v 'Di+86*Tc+50ps' 1.2v 'Di+87*Tc' 1.2v 'Di+87*Tc+50ps' 1.2v 'Di+88*Tc' 1.2v 'Di+88*Tc+50ps' 1.2v 'Di+89*Tc' 1.2v 'Di+89*Tc+50ps' 1.2v 'Di+90*Tc' 1.2v 'Di+90*Tc+50ps' 0v 'Di+91*Tc' 0v 'Di+91*Tc+50ps' 0v 'Di+92*Tc' 0v 'Di+92*Tc+50ps' 1.2v 'Di+93*Tc' 1.2v 'Di+93*Tc+50ps' 0v 'Di+94*Tc' 0v 'Di+94*Tc+50ps' 1.2v 'Di+95*Tc' 1.2v 'Di+95*Tc+50ps' 1.2v 'Di+96*Tc' 1.2v 'Di+96*Tc+50ps' 1.2v 'Di+97*Tc' 1.2v 'Di+97*Tc+50ps' 0v 'Di+98*Tc' 0v 'Di+98*Tc+50ps' 0v 'Di+99*Tc' 0v 'Di+99*Tc+50ps' 0v 'Di+100*Tc' 0v 'Di+100*Tc+50ps' 1.2v 'Di+101*Tc' 1.2v 'Di+101*Tc+50ps' 0v 'Di+102*Tc' 0v 'Di+102*Tc+50ps' 0v 'Di+103*Tc' 0v 'Di+103*Tc+50ps' 1.2v 'Di+104*Tc' 1.2v 'Di+104*Tc+50ps' 1.2v 'Di+105*Tc' 1.2v 'Di+105*Tc+50ps' 0v 'Di+106*Tc' 0v 'Di+106*Tc+50ps' 0v 'Di+107*Tc' 0v 'Di+107*Tc+50ps' 0v 'Di+108*Tc' 0v 'Di+108*Tc+50ps' 0v 'Di+109*Tc' 0v 'Di+109*Tc+50ps' 0v 'Di+110*Tc' 0v)

$The following lines are only to get an example of what the output should look like.
vout_ready_out_exp out_ready_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' 0v 'Di+1*Tc' 0v 'Di+1*Tc+50ps' 0v 'Di+2*Tc' 0v 'Di+2*Tc+50ps' 0v 'Di+3*Tc' 0v 'Di+3*Tc+50ps' 0v 'Di+4*Tc' 0v 'Di+4*Tc+50ps' 0v 'Di+5*Tc' 0v 'Di+5*Tc+50ps' 0v 'Di+6*Tc' 0v 'Di+6*Tc+50ps' 0v 'Di+7*Tc' 0v 'Di+7*Tc+50ps' 0v 'Di+8*Tc' 0v 'Di+8*Tc+50ps' 0v 'Di+9*Tc' 0v 'Di+9*Tc+50ps' 0v 'Di+10*Tc' 0v 'Di+10*Tc+50ps' 0v 'Di+11*Tc' 0v 'Di+11*Tc+50ps' 0v 'Di+12*Tc' 0v 'Di+12*Tc+50ps' 1.2v 'Di+13*Tc' 1.2v 'Di+13*Tc+50ps' 0v 'Di+14*Tc' 0v 'Di+14*Tc+50ps' 0v 'Di+15*Tc' 0v 'Di+15*Tc+50ps' 0v 'Di+16*Tc' 0v 'Di+16*Tc+50ps' 0v 'Di+17*Tc' 0v 'Di+17*Tc+50ps' 0v 'Di+18*Tc' 0v 'Di+18*Tc+50ps' 0v 'Di+19*Tc' 0v 'Di+19*Tc+50ps' 0v 'Di+20*Tc' 0v 'Di+20*Tc+50ps' 0v 'Di+21*Tc' 0v 'Di+21*Tc+50ps' 1.2v 'Di+22*Tc' 1.2v 'Di+22*Tc+50ps' 0v 'Di+23*Tc' 0v 'Di+23*Tc+50ps' 0v 'Di+24*Tc' 0v 'Di+24*Tc+50ps' 0v 'Di+25*Tc' 0v 'Di+25*Tc+50ps' 0v 'Di+26*Tc' 0v 'Di+26*Tc+50ps' 0v 'Di+27*Tc' 0v 'Di+27*Tc+50ps' 0v 'Di+28*Tc' 0v 'Di+28*Tc+50ps' 0v 'Di+29*Tc' 0v 'Di+29*Tc+50ps' 0v 'Di+30*Tc' 0v 'Di+30*Tc+50ps' 0v 'Di+31*Tc' 0v 'Di+31*Tc+50ps' 0v 'Di+32*Tc' 0v 'Di+32*Tc+50ps' 1.2v 'Di+33*Tc' 1.2v 'Di+33*Tc+50ps' 0v 'Di+34*Tc' 0v 'Di+34*Tc+50ps' 0v 'Di+35*Tc' 0v 'Di+35*Tc+50ps' 0v 'Di+36*Tc' 0v 'Di+36*Tc+50ps' 0v 'Di+37*Tc' 0v 'Di+37*Tc+50ps' 0v 'Di+38*Tc' 0v 'Di+38*Tc+50ps' 0v 'Di+39*Tc' 0v 'Di+39*Tc+50ps' 0v 'Di+40*Tc' 0v 'Di+40*Tc+50ps' 1.2v 'Di+41*Tc' 1.2v 'Di+41*Tc+50ps' 0v 'Di+42*Tc' 0v 'Di+42*Tc+50ps' 0v 'Di+43*Tc' 0v 'Di+43*Tc+50ps' 0v 'Di+44*Tc' 0v 'Di+44*Tc+50ps' 0v 'Di+45*Tc' 0v 'Di+45*Tc+50ps' 0v 'Di+46*Tc' 0v 'Di+46*Tc+50ps' 0v 'Di+47*Tc' 0v 'Di+47*Tc+50ps' 0v 'Di+48*Tc' 0v 'Di+48*Tc+50ps' 1.2v 'Di+49*Tc' 1.2v 'Di+49*Tc+50ps' 0v 'Di+50*Tc' 0v 'Di+50*Tc+50ps' 0v 'Di+51*Tc' 0v 'Di+51*Tc+50ps' 0v 'Di+52*Tc' 0v 'Di+52*Tc+50ps' 0v 'Di+53*Tc' 0v 'Di+53*Tc+50ps' 0v 'Di+54*Tc' 0v 'Di+54*Tc+50ps' 0v 'Di+55*Tc' 0v 'Di+55*Tc+50ps' 0v 'Di+56*Tc' 0v 'Di+56*Tc+50ps' 1.2v 'Di+57*Tc' 1.2v 'Di+57*Tc+50ps' 0v 'Di+58*Tc' 0v 'Di+58*Tc+50ps' 0v 'Di+59*Tc' 0v 'Di+59*Tc+50ps' 0v 'Di+60*Tc' 0v 'Di+60*Tc+50ps' 0v 'Di+61*Tc' 0v 'Di+61*Tc+50ps' 0v 'Di+62*Tc' 0v 'Di+62*Tc+50ps' 0v 'Di+63*Tc' 0v 'Di+63*Tc+50ps' 0v 'Di+64*Tc' 0v 'Di+64*Tc+50ps' 0v 'Di+65*Tc' 0v 'Di+65*Tc+50ps' 0v 'Di+66*Tc' 0v 'Di+66*Tc+50ps' 0v 'Di+67*Tc' 0v 'Di+67*Tc+50ps' 0v 'Di+68*Tc' 0v 'Di+68*Tc+50ps' 0v 'Di+69*Tc' 0v 'Di+69*Tc+50ps' 0v 'Di+70*Tc' 0v 'Di+70*Tc+50ps' 0v 'Di+71*Tc' 0v 'Di+71*Tc+50ps' 0v 'Di+72*Tc' 0v 'Di+72*Tc+50ps' 0v 'Di+73*Tc' 0v 'Di+73*Tc+50ps' 0v 'Di+74*Tc' 0v 'Di+74*Tc+50ps' 0v 'Di+75*Tc' 0v 'Di+75*Tc+50ps' 0v 'Di+76*Tc' 0v 'Di+76*Tc+50ps' 0v 'Di+77*Tc' 0v 'Di+77*Tc+50ps' 0v 'Di+78*Tc' 0v 'Di+78*Tc+50ps' 0v 'Di+79*Tc' 0v 'Di+79*Tc+50ps' 0v 'Di+80*Tc' 0v 'Di+80*Tc+50ps' 0v 'Di+81*Tc' 0v 'Di+81*Tc+50ps' 0v 'Di+82*Tc' 0v 'Di+82*Tc+50ps' 0v 'Di+83*Tc' 0v 'Di+83*Tc+50ps' 0v 'Di+84*Tc' 0v 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' 0v 'Di+86*Tc' 0v 'Di+86*Tc+50ps' 0v 'Di+87*Tc' 0v 'Di+87*Tc+50ps' 0v 'Di+88*Tc' 0v 'Di+88*Tc+50ps' 0v 'Di+89*Tc' 0v 'Di+89*Tc+50ps' 0v 'Di+90*Tc' 0v 'Di+90*Tc+50ps' 0v 'Di+91*Tc' 0v 'Di+91*Tc+50ps' 0v 'Di+92*Tc' 0v 'Di+92*Tc+50ps' 1.2v 'Di+93*Tc' 1.2v 'Di+93*Tc+50ps' 0v 'Di+94*Tc' 0v 'Di+94*Tc+50ps' 0v 'Di+95*Tc' 0v 'Di+95*Tc+50ps' 0v 'Di+96*Tc' 0v 'Di+96*Tc+50ps' 0v 'Di+97*Tc' 0v 'Di+97*Tc+50ps' 0v 'Di+98*Tc' 0v 'Di+98*Tc+50ps' 0v 'Di+99*Tc' 0v 'Di+99*Tc+50ps' 0v 'Di+100*Tc' 0v 'Di+100*Tc+50ps' 1.2v 'Di+101*Tc' 1.2v 'Di+101*Tc+50ps' 0v 'Di+102*Tc' 0v 'Di+102*Tc+50ps' 0v 'Di+103*Tc' 0v 'Di+103*Tc+50ps' 0v 'Di+104*Tc' 0v 'Di+104*Tc+50ps' 0v 'Di+105*Tc' 0v 'Di+105*Tc+50ps' 0v 'Di+106*Tc' 0v 'Di+106*Tc+50ps' 0v 'Di+107*Tc' 0v 'Di+107*Tc+50ps' 0v 'Di+108*Tc' 0v 'Di+108*Tc+50ps' 1.2v 'Di+109*Tc' 1.2v 'Di+109*Tc+50ps' 0v 'Di+110*Tc' 0v)

va3_out_exp a3_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' '1.2v/2' 'Di+1*Tc' '1.2v/2' 'Di+1*Tc+50ps' '1.2v/2' 'Di+2*Tc' '1.2v/2' 'Di+2*Tc+50ps' '1.2v/2' 'Di+3*Tc' '1.2v/2' 'Di+3*Tc+50ps' '1.2v/2' 'Di+4*Tc' '1.2v/2' 'Di+4*Tc+50ps' '1.2v/2' 'Di+5*Tc' '1.2v/2' 'Di+5*Tc+50ps' '1.2v/2' 'Di+6*Tc' '1.2v/2' 'Di+6*Tc+50ps' '1.2v/2' 'Di+7*Tc' '1.2v/2' 'Di+7*Tc+50ps' '1.2v/2' 'Di+8*Tc' '1.2v/2' 'Di+8*Tc+50ps' '1.2v/2' 'Di+9*Tc' '1.2v/2' 'Di+9*Tc+50ps' '1.2v/2' 'Di+10*Tc' '1.2v/2' 'Di+10*Tc+50ps' '1.2v/2' 'Di+11*Tc' '1.2v/2' 'Di+11*Tc+50ps' '1.2v/2' 'Di+12*Tc' '1.2v/2' 'Di+12*Tc+50ps' 1.2v 'Di+13*Tc' 1.2v 'Di+13*Tc+50ps' '1.2v/2' 'Di+14*Tc' '1.2v/2' 'Di+14*Tc+50ps' '1.2v/2' 'Di+15*Tc' '1.2v/2' 'Di+15*Tc+50ps' '1.2v/2' 'Di+16*Tc' '1.2v/2' 'Di+16*Tc+50ps' '1.2v/2' 'Di+17*Tc' '1.2v/2' 'Di+17*Tc+50ps' '1.2v/2' 'Di+18*Tc' '1.2v/2' 'Di+18*Tc+50ps' '1.2v/2' 'Di+19*Tc' '1.2v/2' 'Di+19*Tc+50ps' '1.2v/2' 'Di+20*Tc' '1.2v/2' 'Di+20*Tc+50ps' '1.2v/2' 'Di+21*Tc' '1.2v/2' 'Di+21*Tc+50ps' 1.2v 'Di+22*Tc' 1.2v 'Di+22*Tc+50ps' '1.2v/2' 'Di+23*Tc' '1.2v/2' 'Di+23*Tc+50ps' '1.2v/2' 'Di+24*Tc' '1.2v/2' 'Di+24*Tc+50ps' '1.2v/2' 'Di+25*Tc' '1.2v/2' 'Di+25*Tc+50ps' '1.2v/2' 'Di+26*Tc' '1.2v/2' 'Di+26*Tc+50ps' '1.2v/2' 'Di+27*Tc' '1.2v/2' 'Di+27*Tc+50ps' '1.2v/2' 'Di+28*Tc' '1.2v/2' 'Di+28*Tc+50ps' '1.2v/2' 'Di+29*Tc' '1.2v/2' 'Di+29*Tc+50ps' '1.2v/2' 'Di+30*Tc' '1.2v/2' 'Di+30*Tc+50ps' '1.2v/2' 'Di+31*Tc' '1.2v/2' 'Di+31*Tc+50ps' '1.2v/2' 'Di+32*Tc' '1.2v/2' 'Di+32*Tc+50ps' '1.2v/2' 'Di+33*Tc' '1.2v/2' 'Di+33*Tc+50ps' '1.2v/2' 'Di+34*Tc' '1.2v/2' 'Di+34*Tc+50ps' '1.2v/2' 'Di+35*Tc' '1.2v/2' 'Di+35*Tc+50ps' '1.2v/2' 'Di+36*Tc' '1.2v/2' 'Di+36*Tc+50ps' '1.2v/2' 'Di+37*Tc' '1.2v/2' 'Di+37*Tc+50ps' '1.2v/2' 'Di+38*Tc' '1.2v/2' 'Di+38*Tc+50ps' '1.2v/2' 'Di+39*Tc' '1.2v/2' 'Di+39*Tc+50ps' '1.2v/2' 'Di+40*Tc' '1.2v/2' 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' '1.2v/2' 'Di+42*Tc' '1.2v/2' 'Di+42*Tc+50ps' '1.2v/2' 'Di+43*Tc' '1.2v/2' 'Di+43*Tc+50ps' '1.2v/2' 'Di+44*Tc' '1.2v/2' 'Di+44*Tc+50ps' '1.2v/2' 'Di+45*Tc' '1.2v/2' 'Di+45*Tc+50ps' '1.2v/2' 'Di+46*Tc' '1.2v/2' 'Di+46*Tc+50ps' '1.2v/2' 'Di+47*Tc' '1.2v/2' 'Di+47*Tc+50ps' '1.2v/2' 'Di+48*Tc' '1.2v/2' 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' '1.2v/2' 'Di+50*Tc' '1.2v/2' 'Di+50*Tc+50ps' '1.2v/2' 'Di+51*Tc' '1.2v/2' 'Di+51*Tc+50ps' '1.2v/2' 'Di+52*Tc' '1.2v/2' 'Di+52*Tc+50ps' '1.2v/2' 'Di+53*Tc' '1.2v/2' 'Di+53*Tc+50ps' '1.2v/2' 'Di+54*Tc' '1.2v/2' 'Di+54*Tc+50ps' '1.2v/2' 'Di+55*Tc' '1.2v/2' 'Di+55*Tc+50ps' '1.2v/2' 'Di+56*Tc' '1.2v/2' 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' '1.2v/2' 'Di+58*Tc' '1.2v/2' 'Di+58*Tc+50ps' '1.2v/2' 'Di+59*Tc' '1.2v/2' 'Di+59*Tc+50ps' '1.2v/2' 'Di+60*Tc' '1.2v/2' 'Di+60*Tc+50ps' '1.2v/2' 'Di+61*Tc' '1.2v/2' 'Di+61*Tc+50ps' '1.2v/2' 'Di+62*Tc' '1.2v/2' 'Di+62*Tc+50ps' '1.2v/2' 'Di+63*Tc' '1.2v/2' 'Di+63*Tc+50ps' '1.2v/2' 'Di+64*Tc' '1.2v/2' 'Di+64*Tc+50ps' '1.2v/2' 'Di+65*Tc' '1.2v/2' 'Di+65*Tc+50ps' '1.2v/2' 'Di+66*Tc' '1.2v/2' 'Di+66*Tc+50ps' '1.2v/2' 'Di+67*Tc' '1.2v/2' 'Di+67*Tc+50ps' '1.2v/2' 'Di+68*Tc' '1.2v/2' 'Di+68*Tc+50ps' '1.2v/2' 'Di+69*Tc' '1.2v/2' 'Di+69*Tc+50ps' '1.2v/2' 'Di+70*Tc' '1.2v/2' 'Di+70*Tc+50ps' '1.2v/2' 'Di+71*Tc' '1.2v/2' 'Di+71*Tc+50ps' '1.2v/2' 'Di+72*Tc' '1.2v/2' 'Di+72*Tc+50ps' '1.2v/2' 'Di+73*Tc' '1.2v/2' 'Di+73*Tc+50ps' '1.2v/2' 'Di+74*Tc' '1.2v/2' 'Di+74*Tc+50ps' '1.2v/2' 'Di+75*Tc' '1.2v/2' 'Di+75*Tc+50ps' '1.2v/2' 'Di+76*Tc' '1.2v/2' 'Di+76*Tc+50ps' '1.2v/2' 'Di+77*Tc' '1.2v/2' 'Di+77*Tc+50ps' '1.2v/2' 'Di+78*Tc' '1.2v/2' 'Di+78*Tc+50ps' '1.2v/2' 'Di+79*Tc' '1.2v/2' 'Di+79*Tc+50ps' '1.2v/2' 'Di+80*Tc' '1.2v/2' 'Di+80*Tc+50ps' '1.2v/2' 'Di+81*Tc' '1.2v/2' 'Di+81*Tc+50ps' '1.2v/2' 'Di+82*Tc' '1.2v/2' 'Di+82*Tc+50ps' '1.2v/2' 'Di+83*Tc' '1.2v/2' 'Di+83*Tc+50ps' '1.2v/2' 'Di+84*Tc' '1.2v/2' 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' '1.2v/2' 'Di+86*Tc' '1.2v/2' 'Di+86*Tc+50ps' '1.2v/2' 'Di+87*Tc' '1.2v/2' 'Di+87*Tc+50ps' '1.2v/2' 'Di+88*Tc' '1.2v/2' 'Di+88*Tc+50ps' '1.2v/2' 'Di+89*Tc' '1.2v/2' 'Di+89*Tc+50ps' '1.2v/2' 'Di+90*Tc' '1.2v/2' 'Di+90*Tc+50ps' '1.2v/2' 'Di+91*Tc' '1.2v/2' 'Di+91*Tc+50ps' '1.2v/2' 'Di+92*Tc' '1.2v/2' 'Di+92*Tc+50ps' '1.2v/2' 'Di+93*Tc' '1.2v/2' 'Di+93*Tc+50ps' '1.2v/2' 'Di+94*Tc' '1.2v/2' 'Di+94*Tc+50ps' '1.2v/2' 'Di+95*Tc' '1.2v/2' 'Di+95*Tc+50ps' '1.2v/2' 'Di+96*Tc' '1.2v/2' 'Di+96*Tc+50ps' '1.2v/2' 'Di+97*Tc' '1.2v/2' 'Di+97*Tc+50ps' '1.2v/2' 'Di+98*Tc' '1.2v/2' 'Di+98*Tc+50ps' '1.2v/2' 'Di+99*Tc' '1.2v/2' 'Di+99*Tc+50ps' '1.2v/2' 'Di+100*Tc' '1.2v/2' 'Di+100*Tc+50ps' 0v 'Di+101*Tc' 0v 'Di+101*Tc+50ps' '1.2v/2' 'Di+102*Tc' '1.2v/2' 'Di+102*Tc+50ps' '1.2v/2' 'Di+103*Tc' '1.2v/2' 'Di+103*Tc+50ps' '1.2v/2' 'Di+104*Tc' '1.2v/2' 'Di+104*Tc+50ps' '1.2v/2' 'Di+105*Tc' '1.2v/2' 'Di+105*Tc+50ps' '1.2v/2' 'Di+106*Tc' '1.2v/2' 'Di+106*Tc+50ps' '1.2v/2' 'Di+107*Tc' '1.2v/2' 'Di+107*Tc+50ps' '1.2v/2' 'Di+108*Tc' '1.2v/2' 'Di+108*Tc+50ps' 1.2v 'Di+109*Tc' 1.2v 'Di+109*Tc+50ps' '1.2v/2' 'Di+110*Tc' '1.2v/2')
va2_out_exp a2_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' '1.2v/2' 'Di+1*Tc' '1.2v/2' 'Di+1*Tc+50ps' '1.2v/2' 'Di+2*Tc' '1.2v/2' 'Di+2*Tc+50ps' '1.2v/2' 'Di+3*Tc' '1.2v/2' 'Di+3*Tc+50ps' '1.2v/2' 'Di+4*Tc' '1.2v/2' 'Di+4*Tc+50ps' '1.2v/2' 'Di+5*Tc' '1.2v/2' 'Di+5*Tc+50ps' '1.2v/2' 'Di+6*Tc' '1.2v/2' 'Di+6*Tc+50ps' '1.2v/2' 'Di+7*Tc' '1.2v/2' 'Di+7*Tc+50ps' '1.2v/2' 'Di+8*Tc' '1.2v/2' 'Di+8*Tc+50ps' '1.2v/2' 'Di+9*Tc' '1.2v/2' 'Di+9*Tc+50ps' '1.2v/2' 'Di+10*Tc' '1.2v/2' 'Di+10*Tc+50ps' '1.2v/2' 'Di+11*Tc' '1.2v/2' 'Di+11*Tc+50ps' '1.2v/2' 'Di+12*Tc' '1.2v/2' 'Di+12*Tc+50ps' 0v 'Di+13*Tc' 0v 'Di+13*Tc+50ps' '1.2v/2' 'Di+14*Tc' '1.2v/2' 'Di+14*Tc+50ps' '1.2v/2' 'Di+15*Tc' '1.2v/2' 'Di+15*Tc+50ps' '1.2v/2' 'Di+16*Tc' '1.2v/2' 'Di+16*Tc+50ps' '1.2v/2' 'Di+17*Tc' '1.2v/2' 'Di+17*Tc+50ps' '1.2v/2' 'Di+18*Tc' '1.2v/2' 'Di+18*Tc+50ps' '1.2v/2' 'Di+19*Tc' '1.2v/2' 'Di+19*Tc+50ps' '1.2v/2' 'Di+20*Tc' '1.2v/2' 'Di+20*Tc+50ps' '1.2v/2' 'Di+21*Tc' '1.2v/2' 'Di+21*Tc+50ps' 0v 'Di+22*Tc' 0v 'Di+22*Tc+50ps' '1.2v/2' 'Di+23*Tc' '1.2v/2' 'Di+23*Tc+50ps' '1.2v/2' 'Di+24*Tc' '1.2v/2' 'Di+24*Tc+50ps' '1.2v/2' 'Di+25*Tc' '1.2v/2' 'Di+25*Tc+50ps' '1.2v/2' 'Di+26*Tc' '1.2v/2' 'Di+26*Tc+50ps' '1.2v/2' 'Di+27*Tc' '1.2v/2' 'Di+27*Tc+50ps' '1.2v/2' 'Di+28*Tc' '1.2v/2' 'Di+28*Tc+50ps' '1.2v/2' 'Di+29*Tc' '1.2v/2' 'Di+29*Tc+50ps' '1.2v/2' 'Di+30*Tc' '1.2v/2' 'Di+30*Tc+50ps' '1.2v/2' 'Di+31*Tc' '1.2v/2' 'Di+31*Tc+50ps' '1.2v/2' 'Di+32*Tc' '1.2v/2' 'Di+32*Tc+50ps' '1.2v/2' 'Di+33*Tc' '1.2v/2' 'Di+33*Tc+50ps' '1.2v/2' 'Di+34*Tc' '1.2v/2' 'Di+34*Tc+50ps' '1.2v/2' 'Di+35*Tc' '1.2v/2' 'Di+35*Tc+50ps' '1.2v/2' 'Di+36*Tc' '1.2v/2' 'Di+36*Tc+50ps' '1.2v/2' 'Di+37*Tc' '1.2v/2' 'Di+37*Tc+50ps' '1.2v/2' 'Di+38*Tc' '1.2v/2' 'Di+38*Tc+50ps' '1.2v/2' 'Di+39*Tc' '1.2v/2' 'Di+39*Tc+50ps' '1.2v/2' 'Di+40*Tc' '1.2v/2' 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' '1.2v/2' 'Di+42*Tc' '1.2v/2' 'Di+42*Tc+50ps' '1.2v/2' 'Di+43*Tc' '1.2v/2' 'Di+43*Tc+50ps' '1.2v/2' 'Di+44*Tc' '1.2v/2' 'Di+44*Tc+50ps' '1.2v/2' 'Di+45*Tc' '1.2v/2' 'Di+45*Tc+50ps' '1.2v/2' 'Di+46*Tc' '1.2v/2' 'Di+46*Tc+50ps' '1.2v/2' 'Di+47*Tc' '1.2v/2' 'Di+47*Tc+50ps' '1.2v/2' 'Di+48*Tc' '1.2v/2' 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' '1.2v/2' 'Di+50*Tc' '1.2v/2' 'Di+50*Tc+50ps' '1.2v/2' 'Di+51*Tc' '1.2v/2' 'Di+51*Tc+50ps' '1.2v/2' 'Di+52*Tc' '1.2v/2' 'Di+52*Tc+50ps' '1.2v/2' 'Di+53*Tc' '1.2v/2' 'Di+53*Tc+50ps' '1.2v/2' 'Di+54*Tc' '1.2v/2' 'Di+54*Tc+50ps' '1.2v/2' 'Di+55*Tc' '1.2v/2' 'Di+55*Tc+50ps' '1.2v/2' 'Di+56*Tc' '1.2v/2' 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' '1.2v/2' 'Di+58*Tc' '1.2v/2' 'Di+58*Tc+50ps' '1.2v/2' 'Di+59*Tc' '1.2v/2' 'Di+59*Tc+50ps' '1.2v/2' 'Di+60*Tc' '1.2v/2' 'Di+60*Tc+50ps' '1.2v/2' 'Di+61*Tc' '1.2v/2' 'Di+61*Tc+50ps' '1.2v/2' 'Di+62*Tc' '1.2v/2' 'Di+62*Tc+50ps' '1.2v/2' 'Di+63*Tc' '1.2v/2' 'Di+63*Tc+50ps' '1.2v/2' 'Di+64*Tc' '1.2v/2' 'Di+64*Tc+50ps' '1.2v/2' 'Di+65*Tc' '1.2v/2' 'Di+65*Tc+50ps' '1.2v/2' 'Di+66*Tc' '1.2v/2' 'Di+66*Tc+50ps' '1.2v/2' 'Di+67*Tc' '1.2v/2' 'Di+67*Tc+50ps' '1.2v/2' 'Di+68*Tc' '1.2v/2' 'Di+68*Tc+50ps' '1.2v/2' 'Di+69*Tc' '1.2v/2' 'Di+69*Tc+50ps' '1.2v/2' 'Di+70*Tc' '1.2v/2' 'Di+70*Tc+50ps' '1.2v/2' 'Di+71*Tc' '1.2v/2' 'Di+71*Tc+50ps' '1.2v/2' 'Di+72*Tc' '1.2v/2' 'Di+72*Tc+50ps' '1.2v/2' 'Di+73*Tc' '1.2v/2' 'Di+73*Tc+50ps' '1.2v/2' 'Di+74*Tc' '1.2v/2' 'Di+74*Tc+50ps' '1.2v/2' 'Di+75*Tc' '1.2v/2' 'Di+75*Tc+50ps' '1.2v/2' 'Di+76*Tc' '1.2v/2' 'Di+76*Tc+50ps' '1.2v/2' 'Di+77*Tc' '1.2v/2' 'Di+77*Tc+50ps' '1.2v/2' 'Di+78*Tc' '1.2v/2' 'Di+78*Tc+50ps' '1.2v/2' 'Di+79*Tc' '1.2v/2' 'Di+79*Tc+50ps' '1.2v/2' 'Di+80*Tc' '1.2v/2' 'Di+80*Tc+50ps' '1.2v/2' 'Di+81*Tc' '1.2v/2' 'Di+81*Tc+50ps' '1.2v/2' 'Di+82*Tc' '1.2v/2' 'Di+82*Tc+50ps' '1.2v/2' 'Di+83*Tc' '1.2v/2' 'Di+83*Tc+50ps' '1.2v/2' 'Di+84*Tc' '1.2v/2' 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' '1.2v/2' 'Di+86*Tc' '1.2v/2' 'Di+86*Tc+50ps' '1.2v/2' 'Di+87*Tc' '1.2v/2' 'Di+87*Tc+50ps' '1.2v/2' 'Di+88*Tc' '1.2v/2' 'Di+88*Tc+50ps' '1.2v/2' 'Di+89*Tc' '1.2v/2' 'Di+89*Tc+50ps' '1.2v/2' 'Di+90*Tc' '1.2v/2' 'Di+90*Tc+50ps' '1.2v/2' 'Di+91*Tc' '1.2v/2' 'Di+91*Tc+50ps' '1.2v/2' 'Di+92*Tc' '1.2v/2' 'Di+92*Tc+50ps' '1.2v/2' 'Di+93*Tc' '1.2v/2' 'Di+93*Tc+50ps' '1.2v/2' 'Di+94*Tc' '1.2v/2' 'Di+94*Tc+50ps' '1.2v/2' 'Di+95*Tc' '1.2v/2' 'Di+95*Tc+50ps' '1.2v/2' 'Di+96*Tc' '1.2v/2' 'Di+96*Tc+50ps' '1.2v/2' 'Di+97*Tc' '1.2v/2' 'Di+97*Tc+50ps' '1.2v/2' 'Di+98*Tc' '1.2v/2' 'Di+98*Tc+50ps' '1.2v/2' 'Di+99*Tc' '1.2v/2' 'Di+99*Tc+50ps' '1.2v/2' 'Di+100*Tc' '1.2v/2' 'Di+100*Tc+50ps' 1.2v 'Di+101*Tc' 1.2v 'Di+101*Tc+50ps' '1.2v/2' 'Di+102*Tc' '1.2v/2' 'Di+102*Tc+50ps' '1.2v/2' 'Di+103*Tc' '1.2v/2' 'Di+103*Tc+50ps' '1.2v/2' 'Di+104*Tc' '1.2v/2' 'Di+104*Tc+50ps' '1.2v/2' 'Di+105*Tc' '1.2v/2' 'Di+105*Tc+50ps' '1.2v/2' 'Di+106*Tc' '1.2v/2' 'Di+106*Tc+50ps' '1.2v/2' 'Di+107*Tc' '1.2v/2' 'Di+107*Tc+50ps' '1.2v/2' 'Di+108*Tc' '1.2v/2' 'Di+108*Tc+50ps' 1.2v 'Di+109*Tc' 1.2v 'Di+109*Tc+50ps' '1.2v/2' 'Di+110*Tc' '1.2v/2')
va1_out_exp a1_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' '1.2v/2' 'Di+1*Tc' '1.2v/2' 'Di+1*Tc+50ps' '1.2v/2' 'Di+2*Tc' '1.2v/2' 'Di+2*Tc+50ps' '1.2v/2' 'Di+3*Tc' '1.2v/2' 'Di+3*Tc+50ps' '1.2v/2' 'Di+4*Tc' '1.2v/2' 'Di+4*Tc+50ps' '1.2v/2' 'Di+5*Tc' '1.2v/2' 'Di+5*Tc+50ps' '1.2v/2' 'Di+6*Tc' '1.2v/2' 'Di+6*Tc+50ps' '1.2v/2' 'Di+7*Tc' '1.2v/2' 'Di+7*Tc+50ps' '1.2v/2' 'Di+8*Tc' '1.2v/2' 'Di+8*Tc+50ps' '1.2v/2' 'Di+9*Tc' '1.2v/2' 'Di+9*Tc+50ps' '1.2v/2' 'Di+10*Tc' '1.2v/2' 'Di+10*Tc+50ps' '1.2v/2' 'Di+11*Tc' '1.2v/2' 'Di+11*Tc+50ps' '1.2v/2' 'Di+12*Tc' '1.2v/2' 'Di+12*Tc+50ps' 1.2v 'Di+13*Tc' 1.2v 'Di+13*Tc+50ps' '1.2v/2' 'Di+14*Tc' '1.2v/2' 'Di+14*Tc+50ps' '1.2v/2' 'Di+15*Tc' '1.2v/2' 'Di+15*Tc+50ps' '1.2v/2' 'Di+16*Tc' '1.2v/2' 'Di+16*Tc+50ps' '1.2v/2' 'Di+17*Tc' '1.2v/2' 'Di+17*Tc+50ps' '1.2v/2' 'Di+18*Tc' '1.2v/2' 'Di+18*Tc+50ps' '1.2v/2' 'Di+19*Tc' '1.2v/2' 'Di+19*Tc+50ps' '1.2v/2' 'Di+20*Tc' '1.2v/2' 'Di+20*Tc+50ps' '1.2v/2' 'Di+21*Tc' '1.2v/2' 'Di+21*Tc+50ps' 1.2v 'Di+22*Tc' 1.2v 'Di+22*Tc+50ps' '1.2v/2' 'Di+23*Tc' '1.2v/2' 'Di+23*Tc+50ps' '1.2v/2' 'Di+24*Tc' '1.2v/2' 'Di+24*Tc+50ps' '1.2v/2' 'Di+25*Tc' '1.2v/2' 'Di+25*Tc+50ps' '1.2v/2' 'Di+26*Tc' '1.2v/2' 'Di+26*Tc+50ps' '1.2v/2' 'Di+27*Tc' '1.2v/2' 'Di+27*Tc+50ps' '1.2v/2' 'Di+28*Tc' '1.2v/2' 'Di+28*Tc+50ps' '1.2v/2' 'Di+29*Tc' '1.2v/2' 'Di+29*Tc+50ps' '1.2v/2' 'Di+30*Tc' '1.2v/2' 'Di+30*Tc+50ps' '1.2v/2' 'Di+31*Tc' '1.2v/2' 'Di+31*Tc+50ps' '1.2v/2' 'Di+32*Tc' '1.2v/2' 'Di+32*Tc+50ps' '1.2v/2' 'Di+33*Tc' '1.2v/2' 'Di+33*Tc+50ps' '1.2v/2' 'Di+34*Tc' '1.2v/2' 'Di+34*Tc+50ps' '1.2v/2' 'Di+35*Tc' '1.2v/2' 'Di+35*Tc+50ps' '1.2v/2' 'Di+36*Tc' '1.2v/2' 'Di+36*Tc+50ps' '1.2v/2' 'Di+37*Tc' '1.2v/2' 'Di+37*Tc+50ps' '1.2v/2' 'Di+38*Tc' '1.2v/2' 'Di+38*Tc+50ps' '1.2v/2' 'Di+39*Tc' '1.2v/2' 'Di+39*Tc+50ps' '1.2v/2' 'Di+40*Tc' '1.2v/2' 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' '1.2v/2' 'Di+42*Tc' '1.2v/2' 'Di+42*Tc+50ps' '1.2v/2' 'Di+43*Tc' '1.2v/2' 'Di+43*Tc+50ps' '1.2v/2' 'Di+44*Tc' '1.2v/2' 'Di+44*Tc+50ps' '1.2v/2' 'Di+45*Tc' '1.2v/2' 'Di+45*Tc+50ps' '1.2v/2' 'Di+46*Tc' '1.2v/2' 'Di+46*Tc+50ps' '1.2v/2' 'Di+47*Tc' '1.2v/2' 'Di+47*Tc+50ps' '1.2v/2' 'Di+48*Tc' '1.2v/2' 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' '1.2v/2' 'Di+50*Tc' '1.2v/2' 'Di+50*Tc+50ps' '1.2v/2' 'Di+51*Tc' '1.2v/2' 'Di+51*Tc+50ps' '1.2v/2' 'Di+52*Tc' '1.2v/2' 'Di+52*Tc+50ps' '1.2v/2' 'Di+53*Tc' '1.2v/2' 'Di+53*Tc+50ps' '1.2v/2' 'Di+54*Tc' '1.2v/2' 'Di+54*Tc+50ps' '1.2v/2' 'Di+55*Tc' '1.2v/2' 'Di+55*Tc+50ps' '1.2v/2' 'Di+56*Tc' '1.2v/2' 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' '1.2v/2' 'Di+58*Tc' '1.2v/2' 'Di+58*Tc+50ps' '1.2v/2' 'Di+59*Tc' '1.2v/2' 'Di+59*Tc+50ps' '1.2v/2' 'Di+60*Tc' '1.2v/2' 'Di+60*Tc+50ps' '1.2v/2' 'Di+61*Tc' '1.2v/2' 'Di+61*Tc+50ps' '1.2v/2' 'Di+62*Tc' '1.2v/2' 'Di+62*Tc+50ps' '1.2v/2' 'Di+63*Tc' '1.2v/2' 'Di+63*Tc+50ps' '1.2v/2' 'Di+64*Tc' '1.2v/2' 'Di+64*Tc+50ps' '1.2v/2' 'Di+65*Tc' '1.2v/2' 'Di+65*Tc+50ps' '1.2v/2' 'Di+66*Tc' '1.2v/2' 'Di+66*Tc+50ps' '1.2v/2' 'Di+67*Tc' '1.2v/2' 'Di+67*Tc+50ps' '1.2v/2' 'Di+68*Tc' '1.2v/2' 'Di+68*Tc+50ps' '1.2v/2' 'Di+69*Tc' '1.2v/2' 'Di+69*Tc+50ps' '1.2v/2' 'Di+70*Tc' '1.2v/2' 'Di+70*Tc+50ps' '1.2v/2' 'Di+71*Tc' '1.2v/2' 'Di+71*Tc+50ps' '1.2v/2' 'Di+72*Tc' '1.2v/2' 'Di+72*Tc+50ps' '1.2v/2' 'Di+73*Tc' '1.2v/2' 'Di+73*Tc+50ps' '1.2v/2' 'Di+74*Tc' '1.2v/2' 'Di+74*Tc+50ps' '1.2v/2' 'Di+75*Tc' '1.2v/2' 'Di+75*Tc+50ps' '1.2v/2' 'Di+76*Tc' '1.2v/2' 'Di+76*Tc+50ps' '1.2v/2' 'Di+77*Tc' '1.2v/2' 'Di+77*Tc+50ps' '1.2v/2' 'Di+78*Tc' '1.2v/2' 'Di+78*Tc+50ps' '1.2v/2' 'Di+79*Tc' '1.2v/2' 'Di+79*Tc+50ps' '1.2v/2' 'Di+80*Tc' '1.2v/2' 'Di+80*Tc+50ps' '1.2v/2' 'Di+81*Tc' '1.2v/2' 'Di+81*Tc+50ps' '1.2v/2' 'Di+82*Tc' '1.2v/2' 'Di+82*Tc+50ps' '1.2v/2' 'Di+83*Tc' '1.2v/2' 'Di+83*Tc+50ps' '1.2v/2' 'Di+84*Tc' '1.2v/2' 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' '1.2v/2' 'Di+86*Tc' '1.2v/2' 'Di+86*Tc+50ps' '1.2v/2' 'Di+87*Tc' '1.2v/2' 'Di+87*Tc+50ps' '1.2v/2' 'Di+88*Tc' '1.2v/2' 'Di+88*Tc+50ps' '1.2v/2' 'Di+89*Tc' '1.2v/2' 'Di+89*Tc+50ps' '1.2v/2' 'Di+90*Tc' '1.2v/2' 'Di+90*Tc+50ps' '1.2v/2' 'Di+91*Tc' '1.2v/2' 'Di+91*Tc+50ps' '1.2v/2' 'Di+92*Tc' '1.2v/2' 'Di+92*Tc+50ps' '1.2v/2' 'Di+93*Tc' '1.2v/2' 'Di+93*Tc+50ps' '1.2v/2' 'Di+94*Tc' '1.2v/2' 'Di+94*Tc+50ps' '1.2v/2' 'Di+95*Tc' '1.2v/2' 'Di+95*Tc+50ps' '1.2v/2' 'Di+96*Tc' '1.2v/2' 'Di+96*Tc+50ps' '1.2v/2' 'Di+97*Tc' '1.2v/2' 'Di+97*Tc+50ps' '1.2v/2' 'Di+98*Tc' '1.2v/2' 'Di+98*Tc+50ps' '1.2v/2' 'Di+99*Tc' '1.2v/2' 'Di+99*Tc+50ps' '1.2v/2' 'Di+100*Tc' '1.2v/2' 'Di+100*Tc+50ps' 1.2v 'Di+101*Tc' 1.2v 'Di+101*Tc+50ps' '1.2v/2' 'Di+102*Tc' '1.2v/2' 'Di+102*Tc+50ps' '1.2v/2' 'Di+103*Tc' '1.2v/2' 'Di+103*Tc+50ps' '1.2v/2' 'Di+104*Tc' '1.2v/2' 'Di+104*Tc+50ps' '1.2v/2' 'Di+105*Tc' '1.2v/2' 'Di+105*Tc+50ps' '1.2v/2' 'Di+106*Tc' '1.2v/2' 'Di+106*Tc+50ps' '1.2v/2' 'Di+107*Tc' '1.2v/2' 'Di+107*Tc+50ps' '1.2v/2' 'Di+108*Tc' '1.2v/2' 'Di+108*Tc+50ps' 0v 'Di+109*Tc' 0v 'Di+109*Tc+50ps' '1.2v/2' 'Di+110*Tc' '1.2v/2')
va0_out_exp a0_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' '1.2v/2' 'Di+1*Tc' '1.2v/2' 'Di+1*Tc+50ps' '1.2v/2' 'Di+2*Tc' '1.2v/2' 'Di+2*Tc+50ps' '1.2v/2' 'Di+3*Tc' '1.2v/2' 'Di+3*Tc+50ps' '1.2v/2' 'Di+4*Tc' '1.2v/2' 'Di+4*Tc+50ps' '1.2v/2' 'Di+5*Tc' '1.2v/2' 'Di+5*Tc+50ps' '1.2v/2' 'Di+6*Tc' '1.2v/2' 'Di+6*Tc+50ps' '1.2v/2' 'Di+7*Tc' '1.2v/2' 'Di+7*Tc+50ps' '1.2v/2' 'Di+8*Tc' '1.2v/2' 'Di+8*Tc+50ps' '1.2v/2' 'Di+9*Tc' '1.2v/2' 'Di+9*Tc+50ps' '1.2v/2' 'Di+10*Tc' '1.2v/2' 'Di+10*Tc+50ps' '1.2v/2' 'Di+11*Tc' '1.2v/2' 'Di+11*Tc+50ps' '1.2v/2' 'Di+12*Tc' '1.2v/2' 'Di+12*Tc+50ps' 1.2v 'Di+13*Tc' 1.2v 'Di+13*Tc+50ps' '1.2v/2' 'Di+14*Tc' '1.2v/2' 'Di+14*Tc+50ps' '1.2v/2' 'Di+15*Tc' '1.2v/2' 'Di+15*Tc+50ps' '1.2v/2' 'Di+16*Tc' '1.2v/2' 'Di+16*Tc+50ps' '1.2v/2' 'Di+17*Tc' '1.2v/2' 'Di+17*Tc+50ps' '1.2v/2' 'Di+18*Tc' '1.2v/2' 'Di+18*Tc+50ps' '1.2v/2' 'Di+19*Tc' '1.2v/2' 'Di+19*Tc+50ps' '1.2v/2' 'Di+20*Tc' '1.2v/2' 'Di+20*Tc+50ps' '1.2v/2' 'Di+21*Tc' '1.2v/2' 'Di+21*Tc+50ps' 1.2v 'Di+22*Tc' 1.2v 'Di+22*Tc+50ps' '1.2v/2' 'Di+23*Tc' '1.2v/2' 'Di+23*Tc+50ps' '1.2v/2' 'Di+24*Tc' '1.2v/2' 'Di+24*Tc+50ps' '1.2v/2' 'Di+25*Tc' '1.2v/2' 'Di+25*Tc+50ps' '1.2v/2' 'Di+26*Tc' '1.2v/2' 'Di+26*Tc+50ps' '1.2v/2' 'Di+27*Tc' '1.2v/2' 'Di+27*Tc+50ps' '1.2v/2' 'Di+28*Tc' '1.2v/2' 'Di+28*Tc+50ps' '1.2v/2' 'Di+29*Tc' '1.2v/2' 'Di+29*Tc+50ps' '1.2v/2' 'Di+30*Tc' '1.2v/2' 'Di+30*Tc+50ps' '1.2v/2' 'Di+31*Tc' '1.2v/2' 'Di+31*Tc+50ps' '1.2v/2' 'Di+32*Tc' '1.2v/2' 'Di+32*Tc+50ps' '1.2v/2' 'Di+33*Tc' '1.2v/2' 'Di+33*Tc+50ps' '1.2v/2' 'Di+34*Tc' '1.2v/2' 'Di+34*Tc+50ps' '1.2v/2' 'Di+35*Tc' '1.2v/2' 'Di+35*Tc+50ps' '1.2v/2' 'Di+36*Tc' '1.2v/2' 'Di+36*Tc+50ps' '1.2v/2' 'Di+37*Tc' '1.2v/2' 'Di+37*Tc+50ps' '1.2v/2' 'Di+38*Tc' '1.2v/2' 'Di+38*Tc+50ps' '1.2v/2' 'Di+39*Tc' '1.2v/2' 'Di+39*Tc+50ps' '1.2v/2' 'Di+40*Tc' '1.2v/2' 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' '1.2v/2' 'Di+42*Tc' '1.2v/2' 'Di+42*Tc+50ps' '1.2v/2' 'Di+43*Tc' '1.2v/2' 'Di+43*Tc+50ps' '1.2v/2' 'Di+44*Tc' '1.2v/2' 'Di+44*Tc+50ps' '1.2v/2' 'Di+45*Tc' '1.2v/2' 'Di+45*Tc+50ps' '1.2v/2' 'Di+46*Tc' '1.2v/2' 'Di+46*Tc+50ps' '1.2v/2' 'Di+47*Tc' '1.2v/2' 'Di+47*Tc+50ps' '1.2v/2' 'Di+48*Tc' '1.2v/2' 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' '1.2v/2' 'Di+50*Tc' '1.2v/2' 'Di+50*Tc+50ps' '1.2v/2' 'Di+51*Tc' '1.2v/2' 'Di+51*Tc+50ps' '1.2v/2' 'Di+52*Tc' '1.2v/2' 'Di+52*Tc+50ps' '1.2v/2' 'Di+53*Tc' '1.2v/2' 'Di+53*Tc+50ps' '1.2v/2' 'Di+54*Tc' '1.2v/2' 'Di+54*Tc+50ps' '1.2v/2' 'Di+55*Tc' '1.2v/2' 'Di+55*Tc+50ps' '1.2v/2' 'Di+56*Tc' '1.2v/2' 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' '1.2v/2' 'Di+58*Tc' '1.2v/2' 'Di+58*Tc+50ps' '1.2v/2' 'Di+59*Tc' '1.2v/2' 'Di+59*Tc+50ps' '1.2v/2' 'Di+60*Tc' '1.2v/2' 'Di+60*Tc+50ps' '1.2v/2' 'Di+61*Tc' '1.2v/2' 'Di+61*Tc+50ps' '1.2v/2' 'Di+62*Tc' '1.2v/2' 'Di+62*Tc+50ps' '1.2v/2' 'Di+63*Tc' '1.2v/2' 'Di+63*Tc+50ps' '1.2v/2' 'Di+64*Tc' '1.2v/2' 'Di+64*Tc+50ps' '1.2v/2' 'Di+65*Tc' '1.2v/2' 'Di+65*Tc+50ps' '1.2v/2' 'Di+66*Tc' '1.2v/2' 'Di+66*Tc+50ps' '1.2v/2' 'Di+67*Tc' '1.2v/2' 'Di+67*Tc+50ps' '1.2v/2' 'Di+68*Tc' '1.2v/2' 'Di+68*Tc+50ps' '1.2v/2' 'Di+69*Tc' '1.2v/2' 'Di+69*Tc+50ps' '1.2v/2' 'Di+70*Tc' '1.2v/2' 'Di+70*Tc+50ps' '1.2v/2' 'Di+71*Tc' '1.2v/2' 'Di+71*Tc+50ps' '1.2v/2' 'Di+72*Tc' '1.2v/2' 'Di+72*Tc+50ps' '1.2v/2' 'Di+73*Tc' '1.2v/2' 'Di+73*Tc+50ps' '1.2v/2' 'Di+74*Tc' '1.2v/2' 'Di+74*Tc+50ps' '1.2v/2' 'Di+75*Tc' '1.2v/2' 'Di+75*Tc+50ps' '1.2v/2' 'Di+76*Tc' '1.2v/2' 'Di+76*Tc+50ps' '1.2v/2' 'Di+77*Tc' '1.2v/2' 'Di+77*Tc+50ps' '1.2v/2' 'Di+78*Tc' '1.2v/2' 'Di+78*Tc+50ps' '1.2v/2' 'Di+79*Tc' '1.2v/2' 'Di+79*Tc+50ps' '1.2v/2' 'Di+80*Tc' '1.2v/2' 'Di+80*Tc+50ps' '1.2v/2' 'Di+81*Tc' '1.2v/2' 'Di+81*Tc+50ps' '1.2v/2' 'Di+82*Tc' '1.2v/2' 'Di+82*Tc+50ps' '1.2v/2' 'Di+83*Tc' '1.2v/2' 'Di+83*Tc+50ps' '1.2v/2' 'Di+84*Tc' '1.2v/2' 'Di+84*Tc+50ps' 1.2v 'Di+85*Tc' 1.2v 'Di+85*Tc+50ps' '1.2v/2' 'Di+86*Tc' '1.2v/2' 'Di+86*Tc+50ps' '1.2v/2' 'Di+87*Tc' '1.2v/2' 'Di+87*Tc+50ps' '1.2v/2' 'Di+88*Tc' '1.2v/2' 'Di+88*Tc+50ps' '1.2v/2' 'Di+89*Tc' '1.2v/2' 'Di+89*Tc+50ps' '1.2v/2' 'Di+90*Tc' '1.2v/2' 'Di+90*Tc+50ps' '1.2v/2' 'Di+91*Tc' '1.2v/2' 'Di+91*Tc+50ps' '1.2v/2' 'Di+92*Tc' '1.2v/2' 'Di+92*Tc+50ps' '1.2v/2' 'Di+93*Tc' '1.2v/2' 'Di+93*Tc+50ps' '1.2v/2' 'Di+94*Tc' '1.2v/2' 'Di+94*Tc+50ps' '1.2v/2' 'Di+95*Tc' '1.2v/2' 'Di+95*Tc+50ps' '1.2v/2' 'Di+96*Tc' '1.2v/2' 'Di+96*Tc+50ps' '1.2v/2' 'Di+97*Tc' '1.2v/2' 'Di+97*Tc+50ps' '1.2v/2' 'Di+98*Tc' '1.2v/2' 'Di+98*Tc+50ps' '1.2v/2' 'Di+99*Tc' '1.2v/2' 'Di+99*Tc+50ps' '1.2v/2' 'Di+100*Tc' '1.2v/2' 'Di+100*Tc+50ps' 1.2v 'Di+101*Tc' 1.2v 'Di+101*Tc+50ps' '1.2v/2' 'Di+102*Tc' '1.2v/2' 'Di+102*Tc+50ps' '1.2v/2' 'Di+103*Tc' '1.2v/2' 'Di+103*Tc+50ps' '1.2v/2' 'Di+104*Tc' '1.2v/2' 'Di+104*Tc+50ps' '1.2v/2' 'Di+105*Tc' '1.2v/2' 'Di+105*Tc+50ps' '1.2v/2' 'Di+106*Tc' '1.2v/2' 'Di+106*Tc+50ps' '1.2v/2' 'Di+107*Tc' '1.2v/2' 'Di+107*Tc+50ps' '1.2v/2' 'Di+108*Tc' '1.2v/2' 'Di+108*Tc+50ps' 1.2v 'Di+109*Tc' 1.2v 'Di+109*Tc+50ps' '1.2v/2' 'Di+110*Tc' '1.2v/2')

verr_out_exp err_out_exp GND! PWL(0ps 0v Di 0v 'Di+0*Tc+50ps' '1.2v/2' 'Di+1*Tc' '1.2v/2' 'Di+1*Tc+50ps' '1.2v/2' 'Di+2*Tc' '1.2v/2' 'Di+2*Tc+50ps' '1.2v/2' 'Di+3*Tc' '1.2v/2' 'Di+3*Tc+50ps' '1.2v/2' 'Di+4*Tc' '1.2v/2' 'Di+4*Tc+50ps' '1.2v/2' 'Di+5*Tc' '1.2v/2' 'Di+5*Tc+50ps' '1.2v/2' 'Di+6*Tc' '1.2v/2' 'Di+6*Tc+50ps' '1.2v/2' 'Di+7*Tc' '1.2v/2' 'Di+7*Tc+50ps' '1.2v/2' 'Di+8*Tc' '1.2v/2' 'Di+8*Tc+50ps' '1.2v/2' 'Di+9*Tc' '1.2v/2' 'Di+9*Tc+50ps' '1.2v/2' 'Di+10*Tc' '1.2v/2' 'Di+10*Tc+50ps' '1.2v/2' 'Di+11*Tc' '1.2v/2' 'Di+11*Tc+50ps' '1.2v/2' 'Di+12*Tc' '1.2v/2' 'Di+12*Tc+50ps' 0v 'Di+13*Tc' 0v 'Di+13*Tc+50ps' '1.2v/2' 'Di+14*Tc' '1.2v/2' 'Di+14*Tc+50ps' '1.2v/2' 'Di+15*Tc' '1.2v/2' 'Di+15*Tc+50ps' '1.2v/2' 'Di+16*Tc' '1.2v/2' 'Di+16*Tc+50ps' '1.2v/2' 'Di+17*Tc' '1.2v/2' 'Di+17*Tc+50ps' '1.2v/2' 'Di+18*Tc' '1.2v/2' 'Di+18*Tc+50ps' '1.2v/2' 'Di+19*Tc' '1.2v/2' 'Di+19*Tc+50ps' '1.2v/2' 'Di+20*Tc' '1.2v/2' 'Di+20*Tc+50ps' '1.2v/2' 'Di+21*Tc' '1.2v/2' 'Di+21*Tc+50ps' 0v 'Di+22*Tc' 0v 'Di+22*Tc+50ps' '1.2v/2' 'Di+23*Tc' '1.2v/2' 'Di+23*Tc+50ps' '1.2v/2' 'Di+24*Tc' '1.2v/2' 'Di+24*Tc+50ps' '1.2v/2' 'Di+25*Tc' '1.2v/2' 'Di+25*Tc+50ps' '1.2v/2' 'Di+26*Tc' '1.2v/2' 'Di+26*Tc+50ps' '1.2v/2' 'Di+27*Tc' '1.2v/2' 'Di+27*Tc+50ps' '1.2v/2' 'Di+28*Tc' '1.2v/2' 'Di+28*Tc+50ps' '1.2v/2' 'Di+29*Tc' '1.2v/2' 'Di+29*Tc+50ps' '1.2v/2' 'Di+30*Tc' '1.2v/2' 'Di+30*Tc+50ps' '1.2v/2' 'Di+31*Tc' '1.2v/2' 'Di+31*Tc+50ps' '1.2v/2' 'Di+32*Tc' '1.2v/2' 'Di+32*Tc+50ps' 1.2v 'Di+33*Tc' 1.2v 'Di+33*Tc+50ps' '1.2v/2' 'Di+34*Tc' '1.2v/2' 'Di+34*Tc+50ps' '1.2v/2' 'Di+35*Tc' '1.2v/2' 'Di+35*Tc+50ps' '1.2v/2' 'Di+36*Tc' '1.2v/2' 'Di+36*Tc+50ps' '1.2v/2' 'Di+37*Tc' '1.2v/2' 'Di+37*Tc+50ps' '1.2v/2' 'Di+38*Tc' '1.2v/2' 'Di+38*Tc+50ps' '1.2v/2' 'Di+39*Tc' '1.2v/2' 'Di+39*Tc+50ps' '1.2v/2' 'Di+40*Tc' '1.2v/2' 'Di+40*Tc+50ps' 0v 'Di+41*Tc' 0v 'Di+41*Tc+50ps' '1.2v/2' 'Di+42*Tc' '1.2v/2' 'Di+42*Tc+50ps' '1.2v/2' 'Di+43*Tc' '1.2v/2' 'Di+43*Tc+50ps' '1.2v/2' 'Di+44*Tc' '1.2v/2' 'Di+44*Tc+50ps' '1.2v/2' 'Di+45*Tc' '1.2v/2' 'Di+45*Tc+50ps' '1.2v/2' 'Di+46*Tc' '1.2v/2' 'Di+46*Tc+50ps' '1.2v/2' 'Di+47*Tc' '1.2v/2' 'Di+47*Tc+50ps' '1.2v/2' 'Di+48*Tc' '1.2v/2' 'Di+48*Tc+50ps' 0v 'Di+49*Tc' 0v 'Di+49*Tc+50ps' '1.2v/2' 'Di+50*Tc' '1.2v/2' 'Di+50*Tc+50ps' '1.2v/2' 'Di+51*Tc' '1.2v/2' 'Di+51*Tc+50ps' '1.2v/2' 'Di+52*Tc' '1.2v/2' 'Di+52*Tc+50ps' '1.2v/2' 'Di+53*Tc' '1.2v/2' 'Di+53*Tc+50ps' '1.2v/2' 'Di+54*Tc' '1.2v/2' 'Di+54*Tc+50ps' '1.2v/2' 'Di+55*Tc' '1.2v/2' 'Di+55*Tc+50ps' '1.2v/2' 'Di+56*Tc' '1.2v/2' 'Di+56*Tc+50ps' 0v 'Di+57*Tc' 0v 'Di+57*Tc+50ps' '1.2v/2' 'Di+58*Tc' '1.2v/2' 'Di+58*Tc+50ps' '1.2v/2' 'Di+59*Tc' '1.2v/2' 'Di+59*Tc+50ps' '1.2v/2' 'Di+60*Tc' '1.2v/2' 'Di+60*Tc+50ps' '1.2v/2' 'Di+61*Tc' '1.2v/2' 'Di+61*Tc+50ps' '1.2v/2' 'Di+62*Tc' '1.2v/2' 'Di+62*Tc+50ps' '1.2v/2' 'Di+63*Tc' '1.2v/2' 'Di+63*Tc+50ps' '1.2v/2' 'Di+64*Tc' '1.2v/2' 'Di+64*Tc+50ps' '1.2v/2' 'Di+65*Tc' '1.2v/2' 'Di+65*Tc+50ps' '1.2v/2' 'Di+66*Tc' '1.2v/2' 'Di+66*Tc+50ps' '1.2v/2' 'Di+67*Tc' '1.2v/2' 'Di+67*Tc+50ps' '1.2v/2' 'Di+68*Tc' '1.2v/2' 'Di+68*Tc+50ps' '1.2v/2' 'Di+69*Tc' '1.2v/2' 'Di+69*Tc+50ps' '1.2v/2' 'Di+70*Tc' '1.2v/2' 'Di+70*Tc+50ps' '1.2v/2' 'Di+71*Tc' '1.2v/2' 'Di+71*Tc+50ps' '1.2v/2' 'Di+72*Tc' '1.2v/2' 'Di+72*Tc+50ps' '1.2v/2' 'Di+73*Tc' '1.2v/2' 'Di+73*Tc+50ps' '1.2v/2' 'Di+74*Tc' '1.2v/2' 'Di+74*Tc+50ps' '1.2v/2' 'Di+75*Tc' '1.2v/2' 'Di+75*Tc+50ps' '1.2v/2' 'Di+76*Tc' '1.2v/2' 'Di+76*Tc+50ps' '1.2v/2' 'Di+77*Tc' '1.2v/2' 'Di+77*Tc+50ps' '1.2v/2' 'Di+78*Tc' '1.2v/2' 'Di+78*Tc+50ps' '1.2v/2' 'Di+79*Tc' '1.2v/2' 'Di+79*Tc+50ps' '1.2v/2' 'Di+80*Tc' '1.2v/2' 'Di+80*Tc+50ps' '1.2v/2' 'Di+81*Tc' '1.2v/2' 'Di+81*Tc+50ps' '1.2v/2' 'Di+82*Tc' '1.2v/2' 'Di+82*Tc+50ps' '1.2v/2' 'Di+83*Tc' '1.2v/2' 'Di+83*Tc+50ps' '1.2v/2' 'Di+84*Tc' '1.2v/2' 'Di+84*Tc+50ps' 0v 'Di+85*Tc' 0v 'Di+85*Tc+50ps' '1.2v/2' 'Di+86*Tc' '1.2v/2' 'Di+86*Tc+50ps' '1.2v/2' 'Di+87*Tc' '1.2v/2' 'Di+87*Tc+50ps' '1.2v/2' 'Di+88*Tc' '1.2v/2' 'Di+88*Tc+50ps' '1.2v/2' 'Di+89*Tc' '1.2v/2' 'Di+89*Tc+50ps' '1.2v/2' 'Di+90*Tc' '1.2v/2' 'Di+90*Tc+50ps' '1.2v/2' 'Di+91*Tc' '1.2v/2' 'Di+91*Tc+50ps' '1.2v/2' 'Di+92*Tc' '1.2v/2' 'Di+92*Tc+50ps' 1.2v 'Di+93*Tc' 1.2v 'Di+93*Tc+50ps' '1.2v/2' 'Di+94*Tc' '1.2v/2' 'Di+94*Tc+50ps' '1.2v/2' 'Di+95*Tc' '1.2v/2' 'Di+95*Tc+50ps' '1.2v/2' 'Di+96*Tc' '1.2v/2' 'Di+96*Tc+50ps' '1.2v/2' 'Di+97*Tc' '1.2v/2' 'Di+97*Tc+50ps' '1.2v/2' 'Di+98*Tc' '1.2v/2' 'Di+98*Tc+50ps' '1.2v/2' 'Di+99*Tc' '1.2v/2' 'Di+99*Tc+50ps' '1.2v/2' 'Di+100*Tc' '1.2v/2' 'Di+100*Tc+50ps' 0v 'Di+101*Tc' 0v 'Di+101*Tc+50ps' '1.2v/2' 'Di+102*Tc' '1.2v/2' 'Di+102*Tc+50ps' '1.2v/2' 'Di+103*Tc' '1.2v/2' 'Di+103*Tc+50ps' '1.2v/2' 'Di+104*Tc' '1.2v/2' 'Di+104*Tc+50ps' '1.2v/2' 'Di+105*Tc' '1.2v/2' 'Di+105*Tc+50ps' '1.2v/2' 'Di+106*Tc' '1.2v/2' 'Di+106*Tc+50ps' '1.2v/2' 'Di+107*Tc' '1.2v/2' 'Di+107*Tc+50ps' '1.2v/2' 'Di+108*Tc' '1.2v/2' 'Di+108*Tc+50ps' 0v 'Di+109*Tc' 0v 'Di+109*Tc+50ps' '1.2v/2' 'Di+110*Tc' '1.2v/2')

.tr 10ps '112*Tc'  $Run for number of input clock cycles plus 2

.end

